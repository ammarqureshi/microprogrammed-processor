----------------------------------------------------------------------------------
--MUX 3 TO 1
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux3to1_16bits is



end mux3to1_16bits;

architecture Behavioral of mux3to1_16bits is

begin


end Behavioral;

