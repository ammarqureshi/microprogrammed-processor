----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity B_input_logic is

port(B: in std_logic;
s0,s1:in std_logic;
Y: out std_logic

);
end B_input_logic;



architecture Behavioral of B_input_logic is
begin


end Behavioral;

