library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity memory is -- use unsigned for memory address

Port ( address : in  std_logic_vector(15 downto 0);
write_data : in std_logic_vector(15 downto 0);
MemWrite: in std_logic;
read_data : out std_logic_vector(15 downto 0);
CLK: in std_logic);
end memory;


architecture Behavioral of memory is
type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);
-- define type, for memory arrays
begin
mem_process: process (CLK)
-- initialize data memory, X denotes hexadecimal number
variable data_mem : mem_array := (
	X"0000", --0
	X"0000", --1
	X"0241",	--2
	X"0482",	--3
	X"06C3",	--4
	X"0904",	--5
	X"0B45",	--6
	X"0D86",	--7
	X"0FE1",	--8
	X"0000",
	X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",--X"0000", 
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000", 
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
	X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",X"0000", X"0000", X"0000",X"0000"
);
variable addr:integer range 0 to 511;
variable address_out: STD_LOGIC_VECTOR(15 downto 0);

begin -- the following type conversion function is in std_logic_arith
addr:=conv_integer(address(8 downto 0));
address_out:=data_mem(addr);

if MemWrite ='1' then
data_mem(addr):= write_data;

else
read_data<=address_out;

end if;
end process;
end Behavioral;